Library IEEE ;
Use ieee.std_logic_1164.all;

entity BinaryDecimalConverter is
	port(
		
	)